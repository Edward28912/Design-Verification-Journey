`include "uvm_macros.svh"
import uvm_pkg::*;
`include "ram_sequence_lib.sv"
`include "ram_environment.sv"

class ram_write_read_test extends uvm_test;
  `uvm_component_utils(ram_write_read_test)

  ram_env env;
  
  function new(string name = "ram_write_read_test", uvm_component parent);
    super.new(name, parent);
  endfunction
  
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = ram_env::type_id::create("env", this);
  endfunction

  virtual task run_phase(uvm_phase phase);
    ram_write_read_sequence write_read_seq;
    
    phase.raise_objection(this);
    
    #1; env.agent.vif.rstn = 0;
    
    #5; env.agent.vif.rstn = 1;
    `uvm_info(get_type_name(), "Starting write sequence", UVM_MEDIUM)
    
    for(int i = 0; i < 300; i++) begin
      write_read_seq = ram_write_read_sequence::type_id::create("write_read_seq", this);
      write_read_seq.is_random_b = 0;
      write_read_seq.we = 1;
      write_read_seq.addr = i;
      write_read_seq.wdata = i;
      write_read_seq.start(env.agent.sequencer);
    end
    
    for(int i = 0; i < 1300; i++) begin
      write_read_seq = ram_write_read_sequence::type_id::create("write_read_seq", this);
      write_read_seq.is_random_b = 0;
      write_read_seq.we = 0;
      write_read_seq.addr = i;
      write_read_seq.start(env.agent.sequencer);
    end
    
    phase.drop_objection(this);
  endtask

endclass: ram_test
